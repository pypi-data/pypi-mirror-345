* All corners file
.lib init
.include "design.ngspice"
.endl

.lib typical
.lib "sm141064.ngspice" typical
.endl

.lib ff
.lib "sm141064.ngspice" ff
.endl

.lib ss
.lib "sm141064.ngspice" ss
.endl

.lib fs
.lib "sm141064.ngspice" fs
.endl

.lib sf
.lib "sm141064.ngspice" sf
.endl
